module ha(
    input a,b,
    output s,co
    );
assign {co,s}=a+b;
endmodule
